module main

import json

fn (f mut hello.Foo) add(gay &Hello) ?string {
    mut hello := [1,2,3,4]
}

fn main() {
    mut foo := Foo{}
    println(foo.add(Hello))
}